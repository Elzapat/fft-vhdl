library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity iterative_top is
    port (
        
    );
end entity;

architecture top of iterative_top is
begin
end architucture;
